module ProgramCounter
    import DEF::*;
(
    input  logic clk,
    input  logic rst_n,
    input  word  next_pc,
    output word  current_pc
);
    // TODO
endmodule : ProgramCounter
