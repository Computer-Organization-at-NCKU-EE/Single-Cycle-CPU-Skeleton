module BranchComp
    import DEF::*;
(
    input word operand_1,
    input word operand_2,
    BranchCompControlIntf.BranchCompSide control
);
    // TODO
endmodule
