module ImmExt
    import DEF::*;
(
    input  inst_t inst,
    output word   imm_ext_out
);
    // TODO
endmodule
