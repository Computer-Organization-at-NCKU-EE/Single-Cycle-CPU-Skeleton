module LDFilter
    import DEF::*;
(
    input logic [2:0] func3,
    input word in_data,
    output word out_data
);
    // TODO
endmodule
