module ALU
    import DEF::*;  // import package DEF in module header
(
    input alu_opcode_t alu_op,
    input word operand_1,
    input word operand_2,
    output word alu_out
);
    // TODO
endmodule : ALU
